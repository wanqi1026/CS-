LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY F3 IS
PORT(
     D:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
     I15,I14,I13,I12:OUT STD_LOGIC
    );
END F3;

ARCHITECTURE A OF F3 IS
BEGIN
   I15<=D(3);
   I14<=D(2);
   I13<=D(1);
   I12<=D(0);
END A;

