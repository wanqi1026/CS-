LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDR IS
PORT(
	I7,I6,I5,I4: IN STD_LOGIC;
	CF,ZF,SF,OVF,T4,P1,P2,P3: IN STD_LOGIC;
	SE5,SE4,SE3,SE2,SE1,SE0: OUT STD_LOGIC
	);
END ADDR;

ARCHITECTURE A OF ADDR IS
BEGIN
	SE5 <=NOT ((NOT(SF) AND OVF AND P3 AND T4) OR (SF AND NOT(OVF) AND P3 AND T4));
	SE4 <=NOT (CF AND P2 AND T4);
	SE3 <=NOT (I7 AND P1 AND T4);
	SE2 <=NOT (I6 AND P1 AND T4);
	SE1 <=NOT (I5 AND P1 AND T4);
	SE0 <=NOT (I4 AND P1 AND T4);
END A;
