LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY CONTROM IS
PORT(
	ADDR: IN STD_LOGIC_VECTOR(5 DOWNTO 0);--��ַ
	UA: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);--����΢��ַ
	D: OUT STD_LOGIC_VECTOR(20 DOWNTO 0));--΢����
END CONTROM;

ARCHITECTURE A OF CONTROM IS
	SIGNAL DATAOUT: STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN
	PROCESS(ADDR)
	BEGIN
		CASE ADDR IS
			WHEN "000000"=>DATAOUT<="110100100011111101100000000"; --00H ȡָ
			WHEN "000001"=>DATAOUT<="100010100010111011000000000"; --01H IN
			WHEN "000010"=>DATAOUT<="100010100011111110000000000"; --02H MOV
			WHEN "000011"=>DATAOUT<="101000111101110111000001101"; --03H RM_MOV
			WHEN "000100"=>DATAOUT<="101000000011111111000001110"; --04H MR_MOV
			WHEN "000101"=>DATAOUT<="100010000011111111000000000"; --05H RR_MOV
			WHEN "000110"=>DATAOUT<="100000100011111111010000000"; --06H JA
			WHEN "000111"=>DATAOUT<="100000100011111111001000000"; --07H JL
			WHEN "001000"=>DATAOUT<="010000100011111110000000000"; --08H JMP
			WHEN "001001"=>DATAOUT<="100001100111111111000000000"; --09H CMP
			WHEN "001010"=>DATAOUT<="100011101001111111000000000"; --0AH INC
			WHEN "001011"=>DATAOUT<="100011101101111111000000000"; --0BH DEC
			WHEN "001100"=>DATAOUT<="100000000011011111000000000"; --0CH OUT
			WHEN "001101"=>DATAOUT<="100000000011100111000000000"; --0DH RM_MOV(2)
			WHEN "001110"=>DATAOUT<="100010100011110011000000000"; --0EH MR_MOV(2)
			WHEN "010000"=>DATAOUT<="010000100011111110000000000"; --10H JA(2)
			WHEN "100000"=>DATAOUT<="010000100011111110000000000"; --20H JL(2)
			WHEN  OTHERS=>DATAOUT<="100000100011111111000000000";
		END CASE;
		UA(5 DOWNTO 0)<=DATAOUT(5 DOWNTO 0);
		D(20 DOWNTO 0)<=DATAOUT(26 DOWNTO 6);
	END PROCESS;
END A;

