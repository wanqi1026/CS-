LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MCOMMAND IS
PORT(
	T2,T3,T4: IN STD_LOGIC;
	O: IN STD_LOGIC_VECTOR(20 DOWNTO 0);
	P1,P2,P3,LOAD,LDPC,LDAR,LDIR,LDRI,LDPSW,RS_B,S2,S1,S0,ALU_B,SW_B,LED_B,RD_D,CS_D,RAM_B,CS_I,ADDR_B: OUT STD_LOGIC);
END MCOMMAND;

ARCHITECTURE A OF MCOMMAND IS
	SIGNAL DATAOUT: STD_LOGIC_VECTOR(20 DOWNTO 0);
BEGIN
	PROCESS(T2)
	BEGIN
		IF(T2'EVENT AND T2='1') THEN
			DATAOUT(20 DOWNTO 0)<=O(20 DOWNTO 0);
		END IF;
		
		P3<=DATAOUT(0);
		P2<=DATAOUT(1);
		P1<=DATAOUT(2);
		
		ADDR_B<=DATAOUT(3);
		CS_I<=DATAOUT(4);
		RAM_B<=DATAOUT(5);
		CS_D<=NOT(NOT DATAOUT(6) AND T3);
		RD_D<=NOT(NOT DATAOUT(7) AND (T2 OR T3));
		LED_B<=DATAOUT(8);
		SW_B<=DATAOUT(9);
		ALU_B<=DATAOUT(10);
		
		S0<=DATAOUT(11);
		S1<=DATAOUT(12);
		S2<=DATAOUT(13);
		
		RS_B<=DATAOUT(14);
		
		LDPSW<=DATAOUT(15) AND T4;
		
		LDRI<=DATAOUT(16) AND T4;
		LDIR<=DATAOUT(17) AND T3;
		LDAR<=DATAOUT(18) AND T3;
		LDPC<=DATAOUT(19) AND T4;
		LOAD<=DATAOUT(20);
	END PROCESS;
END A;


